library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity decode is
  port (
    clk, rst : in std_logic;
    mem_rd : in std_logic_vector(31 downto 0);
    rs, rt, rd, shamt : out std_logic_vector(4 downto 0);
    imm : out std_logic_vector(15 downto 0);
    target : out std_logic_vector(25 downto 0);
    -- controller
    opcode, funct : out std_logic_vector(5 downto 0);
    instr_clr : in std_logic
  );
end entity;

architecture behavior of decode is
  component flopr_clr
    port (
      clk, rst, clr: in std_logic;
      a : in std_logic_vector(31 downto 0);
      y : out std_logic_vector(31 downto 0)
        );
  end component;

  signal instr0 : std_logic_vector(31 downto 0);
begin
  reg_instr : flopr_clr port map (
    clk => clk, rst => rst, clr => instr_clr,
    a => mem_rd,
    y => instr0
  );

  -- for controller
  opcode <= instr0(31 downto 26);
  rs <= instr0(25 downto 21);
  rt <= instr0(20 downto 16);
  imm <= instr0(15 downto 0);
  target <= instr0(25 downto 0);
  rd <= instr0(15 downto 11);
  shamt <= instr0(10 downto 6);
  funct <= instr0(5 downto 0);
end architecture;
