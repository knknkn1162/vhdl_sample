library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity controller is
  port (
    clk, rst : in std_logic;
    opcode, funct : in std_logic_vector(5 downto 0);
    -- for memadr
    pc_aluout_s, pc_en : out std_logic;
    -- for memwrite
    mem_we: out std_logic;
    -- for writeback
    instr_en, reg_we : out std_logic;
    memrd_aluout_s : out std_logic; -- for lw or addi
    -- for calc
    alucont : out std_logic_vector(2 downto 0);
    rdt_immext_s : out std_logic
  );
end entity;

architecture behavior of controller is
  type statetype is (
    -- soon after the initialization
    InitS, InitFetchS,
    FetchS, DecodeS, AdrCalcS, MemReadS, RegWritebackS,
    MemWriteS,
    -- ExecuteS, ALUWriteBackS,
    -- BranchS,
    AddiExecuteS, AddiWriteBackS
    -- JumpS
  );
  subtype optype is std_logic_vector(5 downto 0);
  constant OP_LW : optype := "100011";
  constant OP_SW : optype := "101011";
  constant OP_ADDI : optype := "001000";
  constant OP_RTYPE : optype := "000000";

  signal state, nextstate : statetype;
begin
  process(clk, rst) begin
    if rst = '1' then
      state <= InitS;
    elsif rising_edge(clk) then
      state <= nextState;
    end if;
  end process;

  -- State Machine
  process(clk, rst, opcode, funct) begin
    case state is
      when InitS =>
        nextState <= InitFetchS;
      when InitFetchS|FetchS =>
        nextState <= DecodeS;
      when DecodeS =>
        case opcode is
          -- lw or sw
          when OP_LW | OP_SW =>
            nextState <= AdrCalcS;
          --when OP_RTYPE =>
          --  nextState <= ExecuteS;
          when OP_ADDI =>
            nextState <= AddiExecuteS;
          when others =>
            nextState <= FetchS;
        end case;
      when AdrCalcS =>
        case opcode is
          when OP_LW =>
            nextState <= MemReadS;
          when OP_SW =>
            nextState <= MemWriteS;
          when others =>
            nextState <= FetchS;
        end case;
      when AddiExecuteS =>
        nextState <= AddiWriteBackS;
      when MemReadS =>
        nextState <= RegWritebackS;
      -- when final state
      when RegWriteBackS | MemWriteS | AddiWriteBackS =>
        nextState <= FetchS;
      -- if undefined
      when others =>
        nextState <= FetchS;
    end case;
  end process;

  -- for sequential logic
  -- ex) D-flipflop enable signal should be turned on before rising_edge(clk)
  process(state)
    variable pc_en0 : std_logic;
    variable instr_en0 : std_logic;
  begin
    pc_en0 := '0';
    instr_en0 := '0';
    case state is
      when InitS =>
        -- pc_en0 := '0';
      when FetchS|InitFetchS =>
        instr_en0 := '1';
      when DecodeS =>
      when AddiExecuteS =>
      when AdrCalcS =>
        -- do nothing
      when MemReadS =>
        -- do nothing
      when MemWriteS | RegWriteBackS | AddiWritebackS =>
        pc_en0 := '1'; -- for fetchS
      when others =>
        -- do nothing;
    end case;

    pc_en <= pc_en0;
    instr_en <= instr_en0;
  end process;

  -- for combinatorial logic
  process(state)
    -- for memadr
    variable pc_aluout_s0 : std_logic;
    -- for memadr
    variable alucont0 : std_logic_vector(2 downto 0);
    variable rdt_immext_s0 : std_logic;
    -- for regwriteback
    variable memrd_aluout_s0 : std_logic;

    -- write in the end of the clk process
    -- for memwrite
    variable mem_we0: std_logic;
    -- for writeback
    variable reg_we0 : std_logic;
  begin
    pc_aluout_s0 := '0';
    alucont0 := "000";
    rdt_immext_s0 := '0';
    memrd_aluout_s0 := '0';
    reg_we0 := '0';
    mem_we0 := '0';
    case state is
      when InitS =>
        -- do nothing
      when InitFetchS =>
        -- do nothing
      when FetchS =>
        -- for decoding
        -- pc_aluout_s0 := '0';
      when DecodeS =>
        -- reg_we0 := '0';
      when AdrCalcS =>
        alucont0 := "010";
        rdt_immext_s0 := '1';
      when AddiExecuteS =>
        alucont0 := "010";
        rdt_immext_s0 := '1';
      when MemReadS =>
        pc_aluout_s0 := '1';
      when MemWriteS =>
        mem_we0 := '1';
        pc_aluout_s0 := '1';
      when RegWriteBackS =>
        reg_we0 := '1';
        -- memrd_aluout_s := '0';
      when AddiWritebackS =>
        reg_we0 := '1';
        memrd_aluout_s0 := '1';
      when others =>
        -- do nothing
    end case;
    pc_aluout_s <= pc_aluout_s0;
    alucont <= alucont0;
    rdt_immext_s <= rdt_immext_s0;
    memrd_aluout_s <= memrd_aluout_s0;
    mem_we <= mem_we0;
    reg_we <= reg_we0;
  end process;
end architecture;
