library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.state_pkg.ALL;

package controller_pkg is
  subtype optype is std_logic_vector(5 downto 0);
  subtype functtype is std_logic_vector(5 downto 0);

  constant OP_LW : optype := "100011"; -- 0x23
  constant OP_SW : optype := "101011"; -- 0x2B
  constant OP_ADDI : optype := "001000"; -- 0x08
  constant OP_ADDIU : optype := "001001"; -- 0x09
  constant OP_ANDI : optype := "001100"; -- 0x0C
  constant OP_SLTI : optype := "001010"; -- 0x0A

  constant OP_RTYPE : optype := "000000";
  constant OP_BEQ : optype := "000100"; -- 0x04
  constant OP_BNE : optype := "000101"; -- 0x05
  constant OP_J : optype := "000010"; -- 0x02

  constant FUNCT_ADD : functtype := "100000"; -- 0x20
  constant FUNCT_ADDU : functtype := "100001"; -- 0x21
  constant FUNCT_AND : functtype := "100100"; -- 0x24
  constant FUNCT_DIV : functtype := "011010"; -- 0x1A
  constant FUNCT_DIVU : functtype := "011011"; -- 0x1B
  constant FUNCT_JR : functtype := "001000"; -- 0x08
  constant FUNCT_NOR : functtype := "100111"; -- 0x27
  constant FUNCT_XOR : functtype := "100110"; -- 0x26
  constant FUNCT_OR : functtype := "100101"; -- 0x25
  constant FUNCT_SLT : functtype := "101010"; -- 0x2A
  constant FUNCT_SLL : functtype := "000000"; -- 0x00
  constant FUNCT_SRL : functtype := "000010"; -- 0x02
  constant FUNCT_SUB : functtype := "100010"; -- 0x22
  constant FUNCT_SUBU : functtype := "100011"; -- 0x23

  function get_nextstate(state: statetype; decs_op: std_logic_vector(5 downto 0); calcs_op: std_logic_vector(5 downto 0); load : std_logic; ena : std_logic; enb : std_logic; is_branch : std_logic) return statetype;
  function get_pc_en(state : statetype) return std_logic;
  function get_instr_clr(stateA: statetype; stateB: statetype; stateC: statetype; is_branch : std_logic) return std_logic;
  function get_pc4_br4_ja_s(state : statetype; opcode : std_logic_vector(5 downto 0); is_branch : std_logic; is_stall : std_logic) return std_logic_vector;
  function get_mem_we(state : statetype) return std_logic;
  function get_alucont(state : statetype; funct : std_logic_vector(5 downto 0)) return std_logic_vector;
  function get_pc_aluout_s(state: statetype) return std_logic;
  function get_rdt_immext_s(state : statetype) return std_logic;
  function get_ena(state: statetype; calcs_opcode : std_logic_vector(5 downto 0); rs : std_logic_vector(4 downto 0); rt: std_logic_vector(4 downto 0); calcs_rt : std_logic_vector(4 downto 0)) return std_logic;
  function get_enb(state1: statetype; state2 : statetype; calcs_opcode : std_logic_vector(5 downto 0)) return std_logic;
  function get_branch_flag(is_equal : std_logic; opcode : std_logic_vector(5 downto 0)) return std_logic;
end package;

package body controller_pkg is
  function get_branch_flag(is_equal : std_logic; opcode : std_logic_vector(5 downto 0)) return std_logic is
    variable is_branch : std_logic;
  begin
    if opcode = OP_BEQ then
      is_branch := is_equal;
    elsif opcode = OP_BNE then
      is_branch := (not is_equal);
    else
      is_branch := '0';
    end if;
    return is_branch;
  end function;

  function get_enb(state1: statetype; state2 : statetype; calcs_opcode : std_logic_vector(5 downto 0)) return std_logic is
    variable enb : std_logic;
  begin
    enb := '1';
    if state1 = MemReadS or state1 = MemWriteBackS then
      -- AdrCalcS is not the end of the state, so the condition `state = AdrCalcS` must not be added
      if state2 = RtypeCalcS or state2 = AddiCalcS or (state2 = AdrCalcS or calcs_opcode = OP_LW) then
        enb := '0';
      end if;
    end if;
    return enb;
  end function;

  function get_ena(state: statetype; calcs_opcode : std_logic_vector(5 downto 0); rs : std_logic_vector(4 downto 0); rt: std_logic_vector(4 downto 0); calcs_rt : std_logic_vector(4 downto 0)) return std_logic is
    variable ena : std_logic;
  begin
    ena := '1';
    if state = AdrCalcS and calcs_opcode = OP_LW then
      if calcs_rt = rt or calcs_rt = rs then
        ena := '0';
      end if;
    end if;
    return ena;
  end function;

  function get_nextstate(state: statetype; decs_op: std_logic_vector(5 downto 0); calcs_op: std_logic_vector(5 downto 0); load : std_logic; ena : std_logic; enb : std_logic; is_branch : std_logic) return statetype is
    variable nextstate : statetype;
  begin
    case state is
      when Wait4S =>
        nextState := Wait3S;
      when Wait3S =>
        nextState := Wait2S;
      when Wait2S =>
        if ena = '0' or enb = '0' then
          nextState := state;
        else
          nextstate := WaitS;
        end if;
      when InitS =>
          nextstate := LoadS;
      when LoadS =>
        nextState := FetchS;
      when WaitS =>
        if enb = '0' then
          nextState := state;
        else
          nextState := FetchS;
        end if;
      when FetchS =>
        if is_branch = '1' then
          nextstate := Wait2S;
        -- stall
        elsif ena = '0' then
          nextState := FetchS;
        else
          nextstate := DecodeS;
        end if;
      when DecodeS =>
        -- stall
        if ena = '1' and enb = '1' then
          case decs_op is
            -- lw or sw
            when OP_LW | OP_SW =>
              nextState := AdrCalcS;
            when OP_RTYPE =>
              nextState := RtypeCalcS;
            when OP_ADDI =>
              nextState := AddiCalcS;
            when OP_BEQ | OP_BNE | OP_J =>
              nextState := WaitS;
            when others =>
              nextState := UnknownS;
          end case;
        else
          -- stay the same state
          nextState := DecodeS;
        end if;
      when AdrCalcS =>
        if enb = '1' then
          case calcs_op is
            when OP_LW =>
              nextState := MemReadS;
            when OP_SW =>
              nextState := MemWriteBackS;
            when others =>
              nextState := UnknownS;
          end case;
        else
          nextState := state;
        end if;
      -- when final state
      when AddiCalcS | RtypeCalcS =>
        if enb = '1' then
          nextState := FetchS;
        else
          nextState := state;
        end if;
      when MemReadS | MemWriteBackS =>
        nextState := FetchS;
      -- if undefined
      when others =>
        nextState := UnknownS;
    end case;
    return nextstate;
  end function;

  function get_pc_en(state : statetype) return std_logic is
    variable ret : std_logic;
  begin
    case state is
      -- when initialization
      when InitS | LoadS | Wait2S | Wait3S | Wait4S =>
        ret := '0';
      when AddiCalcS | RtypeCalcS | MemReadS | MemWriteBackS | WaitS =>
        ret := '1';
      when others =>
        ret := '0';
    end case;
    return ret;
  end function;

  function get_instr_clr(stateA: statetype; stateB: statetype; stateC: statetype; is_branch : std_logic) return std_logic is
    variable ret : std_logic;
  begin
    if stateA = FetchS or stateB = FetchS or stateC = FetchS then
      ret := is_branch;
    else
      ret := '0';
    end if;
    return ret;
  end function;

  function get_pc4_br4_ja_s(state : statetype; opcode : std_logic_vector(5 downto 0); is_branch : std_logic; is_stall : std_logic) return std_logic_vector is
    variable ret : std_logic_vector(1 downto 0);
  begin
    case state is
      when DecodeS =>
        -- "01" : should be taken "00" : shouldnt be taken
        if is_stall = '1' then
          ret := "00";
        elsif opcode = OP_BEQ or opcode = OP_BNE then
          ret := "0" & is_branch;
        elsif opcode = OP_J then
          ret := "10";
        else
          ret := "00";
        end if;
      when others =>
        -- pc+4
        ret := "00";
    end case;
    return ret;
  end function;

  function get_mem_we(state : statetype) return std_logic is
    -- for memwrite
    variable ret: std_logic;
  begin
    case state is
      when MemWriteBackS =>
        ret := '1';
      when others =>
        -- required : MemReadS
        ret := '0';
    end case;
    return ret;
  end function;

  function get_alucont(state : statetype; funct : std_logic_vector(5 downto 0)) return std_logic_vector is
    variable ret : std_logic_vector(2 downto 0);
  begin
    case state is
      when AdrCalcS =>
        ret := "010";
      when RtypeCalcS =>
        case funct is
          when FUNCT_ADD =>
            ret := "010";
          when FUNCT_AND =>
            ret := "000";
          when FUNCT_SUB =>
            ret := "110";
          when FUNCT_SLT =>
            ret := "111";
          when FUNCT_OR =>
            ret := "001";
          when others =>
            ret := "000";
        end case;
      when AddiCalcS =>
        ret := "010";
      when others =>
        ret := "000";
    end case;
    return ret;
  end function;

  function get_pc_aluout_s(state: statetype) return std_logic is
    variable ret : std_logic;
  begin
    case state is
      when MemReadS | MemWriteBackS =>
        ret := '1';
      when others =>
        -- required : FetchS
        ret := '0';
    end case;
    return ret;
  end function;

  function get_rdt_immext_s(state : statetype) return std_logic is
    variable ret : std_logic;
  begin
    case state is
      when AdrCalcS | AddiCalcS =>
        ret := '1';
      when others =>
        -- required : RtypeCalcS
        ret := '0';
    end case;
    return ret;
  end function;
end package body;
