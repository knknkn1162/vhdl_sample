library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.nn_pkg.ALL;

entity sigmoid is
  port (
    a : in std_logic_vector(ASIZE-1 downto 0);
    z : out std_logic_vector(SIZE-1 downto 0)
  );
end entity;

architecture behavior of sigmoid is
  function conv(a : integer) return natural is
    variable b : natural range 0 to 2**SIZE-1;
  begin
    if a < -1419 then b := 0;
    elsif (a >= -1419 and a < -1240) then b := 1;
    elsif (a >= -1240 and a < -1135) then b := 2;
    elsif (a >= -1135 and a < -1061) then b := 3;
    elsif (a >= -1061 and a < -1002) then b := 4;
    elsif (a >= -1002 and a < -955) then b := 5;
    elsif (a >= -955 and a < -914) then b := 6;
    elsif (a >= -914 and a < -879) then b := 7;
    elsif (a >= -879 and a < -848) then b := 8;
    elsif (a >= -848 and a < -820) then b := 9;
    elsif (a >= -820 and a < -794) then b := 10;
    elsif (a >= -794 and a < -771) then b := 11;
    elsif (a >= -771 and a < -750) then b := 12;
    elsif (a >= -750 and a < -730) then b := 13;
    elsif (a >= -730 and a < -711) then b := 14;
    elsif (a >= -711 and a < -693) then b := 15;
    elsif (a >= -693 and a < -677) then b := 16;
    elsif (a >= -677 and a < -661) then b := 17;
    elsif (a >= -661 and a < -646) then b := 18;
    elsif (a >= -646 and a < -632) then b := 19;
    elsif (a >= -632 and a < -618) then b := 20;
    elsif (a >= -618 and a < -605) then b := 21;
    elsif (a >= -605 and a < -593) then b := 22;
    elsif (a >= -593 and a < -581) then b := 23;
    elsif (a >= -581 and a < -569) then b := 24;
    elsif (a >= -569 and a < -558) then b := 25;
    elsif (a >= -558 and a < -547) then b := 26;
    elsif (a >= -547 and a < -537) then b := 27;
    elsif (a >= -537 and a < -527) then b := 28;
    elsif (a >= -527 and a < -517) then b := 29;
    elsif (a >= -517 and a < -507) then b := 30;
    elsif (a >= -507 and a < -498) then b := 31;
    elsif (a >= -498 and a < -489) then b := 32;
    elsif (a >= -489 and a < -480) then b := 33;
    elsif (a >= -480 and a < -472) then b := 34;
    elsif (a >= -472 and a < -463) then b := 35;
    elsif (a >= -463 and a < -455) then b := 36;
    elsif (a >= -455 and a < -447) then b := 37;
    elsif (a >= -447 and a < -439) then b := 38;
    elsif (a >= -439 and a < -432) then b := 39;
    elsif (a >= -432 and a < -424) then b := 40;
    elsif (a >= -424 and a < -417) then b := 41;
    elsif (a >= -417 and a < -410) then b := 42;
    elsif (a >= -410 and a < -403) then b := 43;
    elsif (a >= -403 and a < -396) then b := 44;
    elsif (a >= -396 and a < -389) then b := 45;
    elsif (a >= -389 and a < -382) then b := 46;
    elsif (a >= -382 and a < -375) then b := 47;
    elsif (a >= -375 and a < -369) then b := 48;
    elsif (a >= -369 and a < -362) then b := 49;
    elsif (a >= -362 and a < -356) then b := 50;
    elsif (a >= -356 and a < -350) then b := 51;
    elsif (a >= -350 and a < -344) then b := 52;
    elsif (a >= -344 and a < -338) then b := 53;
    elsif (a >= -338 and a < -332) then b := 54;
    elsif (a >= -332 and a < -326) then b := 55;
    elsif (a >= -326 and a < -320) then b := 56;
    elsif (a >= -320 and a < -314) then b := 57;
    elsif (a >= -314 and a < -309) then b := 58;
    elsif (a >= -309 and a < -303) then b := 59;
    elsif (a >= -303 and a < -298) then b := 60;
    elsif (a >= -298 and a < -292) then b := 61;
    elsif (a >= -292 and a < -287) then b := 62;
    elsif (a >= -287 and a < -281) then b := 63;
    elsif (a >= -281 and a < -276) then b := 64;
    elsif (a >= -276 and a < -271) then b := 65;
    elsif (a >= -271 and a < -265) then b := 66;
    elsif (a >= -265 and a < -260) then b := 67;
    elsif (a >= -260 and a < -255) then b := 68;
    elsif (a >= -255 and a < -250) then b := 69;
    elsif (a >= -250 and a < -245) then b := 70;
    elsif (a >= -245 and a < -240) then b := 71;
    elsif (a >= -240 and a < -235) then b := 72;
    elsif (a >= -235 and a < -230) then b := 73;
    elsif (a >= -230 and a < -226) then b := 74;
    elsif (a >= -226 and a < -221) then b := 75;
    elsif (a >= -221 and a < -216) then b := 76;
    elsif (a >= -216 and a < -211) then b := 77;
    elsif (a >= -211 and a < -207) then b := 78;
    elsif (a >= -207 and a < -202) then b := 79;
    elsif (a >= -202 and a < -197) then b := 80;
    elsif (a >= -197 and a < -193) then b := 81;
    elsif (a >= -193 and a < -188) then b := 82;
    elsif (a >= -188 and a < -183) then b := 83;
    elsif (a >= -183 and a < -179) then b := 84;
    elsif (a >= -179 and a < -174) then b := 85;
    elsif (a >= -174 and a < -170) then b := 86;
    elsif (a >= -170 and a < -166) then b := 87;
    elsif (a >= -166 and a < -161) then b := 88;
    elsif (a >= -161 and a < -157) then b := 89;
    elsif (a >= -157 and a < -152) then b := 90;
    elsif (a >= -152 and a < -148) then b := 91;
    elsif (a >= -148 and a < -144) then b := 92;
    elsif (a >= -144 and a < -139) then b := 93;
    elsif (a >= -139 and a < -135) then b := 94;
    elsif (a >= -135 and a < -131) then b := 95;
    elsif (a >= -131 and a < -127) then b := 96;
    elsif (a >= -127 and a < -122) then b := 97;
    elsif (a >= -122 and a < -118) then b := 98;
    elsif (a >= -118 and a < -114) then b := 99;
    elsif (a >= -114 and a < -110) then b := 100;
    elsif (a >= -110 and a < -105) then b := 101;
    elsif (a >= -105 and a < -101) then b := 102;
    elsif (a >= -101 and a < -97) then b := 103;
    elsif (a >= -97 and a < -93) then b := 104;
    elsif (a >= -93 and a < -89) then b := 105;
    elsif (a >= -89 and a < -85) then b := 106;
    elsif (a >= -85 and a < -81) then b := 107;
    elsif (a >= -81 and a < -77) then b := 108;
    elsif (a >= -77 and a < -72) then b := 109;
    elsif (a >= -72 and a < -68) then b := 110;
    elsif (a >= -68 and a < -64) then b := 111;
    elsif (a >= -64 and a < -60) then b := 112;
    elsif (a >= -60 and a < -56) then b := 113;
    elsif (a >= -56 and a < -52) then b := 114;
    elsif (a >= -52 and a < -48) then b := 115;
    elsif (a >= -48 and a < -44) then b := 116;
    elsif (a >= -44 and a < -40) then b := 117;
    elsif (a >= -40 and a < -36) then b := 118;
    elsif (a >= -36 and a < -32) then b := 119;
    elsif (a >= -32 and a < -28) then b := 120;
    elsif (a >= -28 and a < -24) then b := 121;
    elsif (a >= -24 and a < -20) then b := 122;
    elsif (a >= -20 and a < -16) then b := 123;
    elsif (a >= -16 and a < -12) then b := 124;
    elsif (a >= -12 and a < -8) then b := 125;
    elsif (a >= -8 and a < -4) then b := 126;
    elsif (a >= -4 and a < 0) then b := 127;
    elsif (a >= 0 and a < 4) then b := 128;
    elsif (a >= 4 and a < 8) then b := 129;
    elsif (a >= 8 and a < 12) then b := 130;
    elsif (a >= 12 and a < 16) then b := 131;
    elsif (a >= 16 and a < 20) then b := 132;
    elsif (a >= 20 and a < 24) then b := 133;
    elsif (a >= 24 and a < 28) then b := 134;
    elsif (a >= 28 and a < 32) then b := 135;
    elsif (a >= 32 and a < 36) then b := 136;
    elsif (a >= 36 and a < 40) then b := 137;
    elsif (a >= 40 and a < 44) then b := 138;
    elsif (a >= 44 and a < 48) then b := 139;
    elsif (a >= 48 and a < 52) then b := 140;
    elsif (a >= 52 and a < 56) then b := 141;
    elsif (a >= 56 and a < 60) then b := 142;
    elsif (a >= 60 and a < 64) then b := 143;
    elsif (a >= 64 and a < 68) then b := 144;
    elsif (a >= 68 and a < 72) then b := 145;
    elsif (a >= 72 and a < 77) then b := 146;
    elsif (a >= 77 and a < 81) then b := 147;
    elsif (a >= 81 and a < 85) then b := 148;
    elsif (a >= 85 and a < 89) then b := 149;
    elsif (a >= 89 and a < 93) then b := 150;
    elsif (a >= 93 and a < 97) then b := 151;
    elsif (a >= 97 and a < 101) then b := 152;
    elsif (a >= 101 and a < 105) then b := 153;
    elsif (a >= 105 and a < 110) then b := 154;
    elsif (a >= 110 and a < 114) then b := 155;
    elsif (a >= 114 and a < 118) then b := 156;
    elsif (a >= 118 and a < 122) then b := 157;
    elsif (a >= 122 and a < 127) then b := 158;
    elsif (a >= 127 and a < 131) then b := 159;
    elsif (a >= 131 and a < 135) then b := 160;
    elsif (a >= 135 and a < 139) then b := 161;
    elsif (a >= 139 and a < 144) then b := 162;
    elsif (a >= 144 and a < 148) then b := 163;
    elsif (a >= 148 and a < 152) then b := 164;
    elsif (a >= 152 and a < 157) then b := 165;
    elsif (a >= 157 and a < 161) then b := 166;
    elsif (a >= 161 and a < 166) then b := 167;
    elsif (a >= 166 and a < 170) then b := 168;
    elsif (a >= 170 and a < 174) then b := 169;
    elsif (a >= 174 and a < 179) then b := 170;
    elsif (a >= 179 and a < 183) then b := 171;
    elsif (a >= 183 and a < 188) then b := 172;
    elsif (a >= 188 and a < 193) then b := 173;
    elsif (a >= 193 and a < 197) then b := 174;
    elsif (a >= 197 and a < 202) then b := 175;
    elsif (a >= 202 and a < 207) then b := 176;
    elsif (a >= 207 and a < 211) then b := 177;
    elsif (a >= 211 and a < 216) then b := 178;
    elsif (a >= 216 and a < 221) then b := 179;
    elsif (a >= 221 and a < 226) then b := 180;
    elsif (a >= 226 and a < 230) then b := 181;
    elsif (a >= 230 and a < 235) then b := 182;
    elsif (a >= 235 and a < 240) then b := 183;
    elsif (a >= 240 and a < 245) then b := 184;
    elsif (a >= 245 and a < 250) then b := 185;
    elsif (a >= 250 and a < 255) then b := 186;
    elsif (a >= 255 and a < 260) then b := 187;
    elsif (a >= 260 and a < 265) then b := 188;
    elsif (a >= 265 and a < 271) then b := 189;
    elsif (a >= 271 and a < 276) then b := 190;
    elsif (a >= 276 and a < 281) then b := 191;
    elsif (a >= 281 and a < 287) then b := 192;
    elsif (a >= 287 and a < 292) then b := 193;
    elsif (a >= 292 and a < 298) then b := 194;
    elsif (a >= 298 and a < 303) then b := 195;
    elsif (a >= 303 and a < 309) then b := 196;
    elsif (a >= 309 and a < 314) then b := 197;
    elsif (a >= 314 and a < 320) then b := 198;
    elsif (a >= 320 and a < 326) then b := 199;
    elsif (a >= 326 and a < 332) then b := 200;
    elsif (a >= 332 and a < 338) then b := 201;
    elsif (a >= 338 and a < 344) then b := 202;
    elsif (a >= 344 and a < 350) then b := 203;
    elsif (a >= 350 and a < 356) then b := 204;
    elsif (a >= 356 and a < 362) then b := 205;
    elsif (a >= 362 and a < 369) then b := 206;
    elsif (a >= 369 and a < 375) then b := 207;
    elsif (a >= 375 and a < 382) then b := 208;
    elsif (a >= 382 and a < 389) then b := 209;
    elsif (a >= 389 and a < 396) then b := 210;
    elsif (a >= 396 and a < 403) then b := 211;
    elsif (a >= 403 and a < 410) then b := 212;
    elsif (a >= 410 and a < 417) then b := 213;
    elsif (a >= 417 and a < 424) then b := 214;
    elsif (a >= 424 and a < 432) then b := 215;
    elsif (a >= 432 and a < 439) then b := 216;
    elsif (a >= 439 and a < 447) then b := 217;
    elsif (a >= 447 and a < 455) then b := 218;
    elsif (a >= 455 and a < 463) then b := 219;
    elsif (a >= 463 and a < 472) then b := 220;
    elsif (a >= 472 and a < 480) then b := 221;
    elsif (a >= 480 and a < 489) then b := 222;
    elsif (a >= 489 and a < 498) then b := 223;
    elsif (a >= 498 and a < 507) then b := 224;
    elsif (a >= 507 and a < 517) then b := 225;
    elsif (a >= 517 and a < 527) then b := 226;
    elsif (a >= 527 and a < 537) then b := 227;
    elsif (a >= 537 and a < 547) then b := 228;
    elsif (a >= 547 and a < 558) then b := 229;
    elsif (a >= 558 and a < 569) then b := 230;
    elsif (a >= 569 and a < 581) then b := 231;
    elsif (a >= 581 and a < 593) then b := 232;
    elsif (a >= 593 and a < 605) then b := 233;
    elsif (a >= 605 and a < 618) then b := 234;
    elsif (a >= 618 and a < 632) then b := 235;
    elsif (a >= 632 and a < 646) then b := 236;
    elsif (a >= 646 and a < 661) then b := 237;
    elsif (a >= 661 and a < 677) then b := 238;
    elsif (a >= 677 and a < 693) then b := 239;
    elsif (a >= 693 and a < 711) then b := 240;
    elsif (a >= 711 and a < 730) then b := 241;
    elsif (a >= 730 and a < 750) then b := 242;
    elsif (a >= 750 and a < 771) then b := 243;
    elsif (a >= 771 and a < 794) then b := 244;
    elsif (a >= 794 and a < 820) then b := 245;
    elsif (a >= 820 and a < 848) then b := 246;
    elsif (a >= 848 and a < 879) then b := 247;
    elsif (a >= 879 and a < 914) then b := 248;
    elsif (a >= 914 and a < 955) then b := 249;
    elsif (a >= 955 and a < 1002) then b := 250;
    elsif (a >= 1002 and a < 1061) then b := 251;
    elsif (a >= 1061 and a < 1135) then b := 252;
    elsif (a >= 1135 and a < 1240) then b := 253;
    elsif (a >= 1240 and a < 1419) then b := 254;
    else b := 255;
  end if;
  return b;
  end function;
begin
  process(a) begin
    if is_X(a) then
      z <= (others => '-');
    else
      z <= std_logic_vector(to_unsigned(conv(to_integer(signed(a))), SIZE));
    end if;
  end process;
end architecture;
